module Image_Processing();



endmodule
